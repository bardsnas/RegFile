module DE1_SoC